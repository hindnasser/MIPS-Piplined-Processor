module ALUcontrol ();

endmodule
