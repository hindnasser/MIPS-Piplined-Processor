module ZeroExtension ();
 
endmodule
