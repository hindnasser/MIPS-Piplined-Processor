module MEM_WB_Register ();
endmodule
