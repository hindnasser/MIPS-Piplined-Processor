module ShiftLift2 ();

endmodule
