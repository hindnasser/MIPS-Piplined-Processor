module AddressAdder ();

endmodule
