module HazardDetectionUnit ();

endmodule
