module ALU (EXE_Result, EXE_Zero, Overflow, Op1, Op2, operation, shamt, clk);

// input
	input [31:0] Op1, Op2;
	input [3:0] operation;
	input [4:0] shamt;
	input clk;
	
// output
	output reg [31:0] EXE_Result;
	output reg EXE_Zero, Overflow;
	
// cases

	always @ (posedge clk) begin
		case (operation)

//			// unsigned addition 
//			4'h0:
//				begin
//					EXE_Result <= Op1 + Op2;
//					EXE_Zero <= 0;
//					Overflow <= 0;
//				end

			// no Operation 
				4'h0:
					begin
						EXE_Result <= 0;
						EXE_Zero <= 0;
						Overflow <= 0;
					end
				
			//shift lift 16 for Op2
			4'h11:
				begin
					EXE_Result <= Op2 << 16;
					EXE_Zero <= 0;
					Overflow <= 0;
				end
				
			//Or 
			4'h3:
				begin
					EXE_Result <= Op1 | Op2;
					EXE_Zero <= 0;
					Overflow <= 0;
				end
				
			//signed addition
			4'h4:
				begin
					EXE_Result <= Op1 + Op2;
					EXE_Zero <= 0;
				   // To detect overflow
					if (Op1[31] == Op2[31] && EXE_Result[31] == Op1[31]) 
							Overflow <= 0;
							
					else Overflow <= 1;
				end
				
			//and 
			4'h5:
				begin
					EXE_Result <= Op1 & Op2;
					EXE_Zero <= 0;
					Overflow <= 0;
				end
				
//			//Unsigned Subtract
//			4'h6:
//				begin
//					EXE_Result <= Op2 - Op1;
//					//to detect the EXE_Zero value
//					if(EXE_Result == 32'h0)
//						EXE_Zero <= 1;
//						
//					else EXE_Zero <= 0;
//					Overflow <= 0;
//				end
				
				
			//Signed Subtract
			4'h7:
				begin
					EXE_Result <= Op2 - Op1;
					
					//to detect overflow
					if(Op2[31] != Op1[31] && EXE_Result[31]== Op1[31])
						Overflow <= 1;
						
					else Overflow <= 0;
					
					//to detect the EXE_Zero bit
					if(EXE_Result == 32'h0 && Overflow == 0)
						EXE_Zero <= 1;
						
					else EXE_Zero <= 0;
				end
				
			//Shift lift 
			4'h8:
				begin
					EXE_Result <= Op2 << shamt;
					EXE_Zero <= 0;
					Overflow <= 0;
				end
			
			//Shift right
			4'h9:
				begin
					EXE_Result <= Op2 >> shamt;
					EXE_Zero <= 0;
					Overflow <=0;
				end
				
			//Set less than
			4'h12:
				begin
					if($signed (Op1) < $signed (Op2)) EXE_Result <= 1;
					else EXE_Result <= 0; 
					EXE_Zero <= 0;
					Overflow <=0;
				end
				
			//Set less than unsigned
			4'h13:
				begin
					if( Op1 < Op2) EXE_Result <= 1;
					else EXE_Result <= 0;
					EXE_Zero <= 0;
					Overflow <=0;
				end
				
			//Nor
			4'h14:
				begin
					EXE_Result <= ~(Op1 | Op2);
					EXE_Zero <= 0;
					Overflow <=0;
				end
				
			//Passing rt for Jr
			4'h15:
				begin
					EXE_Result <= Op2;
					EXE_Zero <= 0;
					Overflow <=0;
				end
							
		endcase
		
	end
		
endmodule
