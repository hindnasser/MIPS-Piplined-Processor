module EXE_MEM_Register ();
endmodule
