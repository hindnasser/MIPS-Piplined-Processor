module PCAdder ();

endmodule
