module SignExtension ();

endmodule
