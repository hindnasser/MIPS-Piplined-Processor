module Top (PC_value);

// input
	input [31:0] PC_value;
   
// clock
	wire clk;
	clock c(clk);
	
// wires
	// IF Stage
	wire [31:0] instruction, PCplus4, program_counter, Mem_BranchAddress, PCSrc;
	wire PC_Src;
	
	//IF_ID_Register
	wire [4:0] IF_ID_Rs, IF_ID_Rt, IF_ID_Rd, IF_ID_Shamt;
	wire [5:0] IF_ID_Func, IF_ID_Opcode;
	wire [15:0] IF_ID_Immediate;
	wire [25:0] IF_ID_Address;
	wire [31:0] IF_ID_PCplus4Out;
	
	// ID Stage
	wire [31:0] SignedImmediate, UnsignedImmediate, ReadData1, ReadData2, ExtendedImm;					
	wire RegDst, RegWrite, MemtoReg, Jump, JmpandLink, MemRead, MemWrite, BranchEqual, BranchnotEqual, ALUop, ALUSrc, floatop, Issigned;
	
	// ID_EXE_Register
	wire ID_EXE_RegDst, ID_EXE_RegWrite, ID_EXE_MemtoReg, ID_EXE_JmpandLink, ID_EXE_MemRead, ID_EXE_MemWrite, ID_EXE_BranchEqual, ID_EXE_BranchnotEqual,
		  ID_EXE_ALUSrc;
	wire [5:0] ID_EXE_Func;
	wire [31:0] ID_EXE_PCplus4, ID_EXE_Rs, ID_EXE_Rt, ID_EXE_ExtendedImm;
	wire [4:0] ID_EXE_Shamt, ID_EXE_Rd; 
	// EXE Stage
	wire [31:0] ALUOut_EXEC, Op2Srcs, Op1, Op2, BranchAdd, EXE_BranchAddress;
	wire EXE_Zero, Overflow, forwardOp1, forwardOp2;
	wire [4:0] EXE_DstReg;
	
	// EXE_MEM_Register
	wire [31:0] EXE_MEM_Result, EXE_MEM_BranchAddress, EXE_MEM_Rt;
	wire EXE_MEM_Zero, EXE_MEM_BranchEqual, EXE_MEM_BranchnotEqual, EXE_MEM_MemRead, EXE_MEM_MemWrite, EXE_MEM_MemtoReg, EXE_MEM_RegWrite; 
	wire [4:0] EXE_MEM_DstReg, EXE_MEM_Rd;
	
	// MEM Stage
	wire [31:0] MEM_Result;
	wire BranchEqualResult, BranchnotEqualResult;
	
	// MEM_ WB_Register
	wire [31:0] MEM_WB_MemData, MEM_WB_ALUData;
	wire [4:0] MEM_WB_Rd, MEM_WB_DstReg;
	wire MEM_WB_MemtoReg, MEM_WB_RegWrite;
	
	// WB Stage
	wire [31:0] WB_Data;
	
// IF Stage
	PC_MUX pcmux (PCSrc, PC_value, Mem_BranchAddress, PC_Src);
	PC_Reg pcreg (program_counter, PCSrc);
	PCAdder pcadd (PCplus4, program_counter);
	instructionMemory imem (instruction, program_counter);

// IF_ID_Register
	IF_ID_Register ifidr (IF_ID_Rs, IF_ID_Rt, IF_ID_Rd, IF_ID_Opcode, IF_ID_Shamt, IF_ID_Func, IF_ID_Immediate,
								 IF_ID_Address, IF_ID_PCplus4Out, instruction, clk, PCplus4); 
	
// ID Stage
	ControlUnit cu (RegDst, RegWrite, MemtoReg, Jump, JmpandLink, MemRead, MemWrite, BranchEqual, BranchnotEqual, ALUop, ALUSrc, floatop, Issigned, IF_ID_Opcode);
	SignExtension se (SignedImmediate, IF_ID_Immediate);
	ZeroExtension ze (UnsignedImmediate, IF_ID_Immediate );
	Ext_MUX extmux (ExtendedImm, SignedImmediate, UnsignedImmediate, Issigned, clk);
	RegisterFile regFile (ReadData1, ReadData2, clk, IF_ID_Rs, IF_ID_Rt, WB_DstReg, WB_Data, RegWrite);//here
	// floating register file
	// Rs_MUX
	// Rs_MUX rsmux (ID_Rs, ReadData1, FPReadData1, floatop, clk);
	// Rt_MUx
	// Rt_MUX rtmux (ID_Rt, ReadData2, FPReadData2, floatop, clk);
	
// ID_EXE_Register
	ID_EXE_Register idexer (ID_EXE_Func, ID_EXE_PCplus4, ID_EXE_Rs, ID_EXE_Rt, ID_EXE_Rd, ID_EXE_ExtendedImm, ID_EXE_Shamt, ID_EXE_RegDst, ID_EXE_RegWrite, 
	                        ID_EXE_MemtoReg, ID_EXE_JmpandLink, ID_EXE_MemRead, ID_EXE_MemWrite, ID_EXE_BranchEqual, ID_EXE_BranchnotEqual, ID_EXE_ALUop, 
									ID_EXE_ALUSrc, IF_ID_Shamt, IF_ID_Func, IF_ID_PCplus4, ReadData1, ReadData2, IF_ID_Rd, ExtendedImm, RegDst, RegWrite, MemtoReg,
									// change ReadData1 and ReadData2 to ID_Rs and ID_Rt after adding floating point registerFile
									JmpandLink, MemRead, MemWrite, BranchEqual, BranchnotEqual, ALUop, ALUSrc, clk);
												
// EXE Stage
	Op2Src_MUX op2srcmux (Op2Src, ID_EXE_Rt, ID_EXE_ExtendedImm, ID_EXE_ALUSrc, clk);
	ForOp1_MUX forop1mux (Op1, ID_EXE_Rs, WB_Data, EXE_MEM_Result, forwardOp1, clk);
	ForOp2_MUX forop2mux (Op2, Op2Src, WB_Data, EXE_MEM_Result, forwardOp2, clk);
	DstReg_MUX dstregmux (EXE_DstReg, ID_EXE_Rt, ID_EXE_Rd, ID_EXE_RegDst, clk);

	AddressAdder addadd (EXE_BranchAddress, ID_EXE_PCplus4, BranchAdd);
	ALU alu (ALUOut_EXEC, EXE_Zero, Overflow, Op1, Op2, 4'h4, ID_EXE_Shamt, clk);//here
	// change nmber to operation after adding the alu control
	ForwardingUnit forunit (forwardOp1, forwardOp2, ID_EXE_Rs, ID_EXE_Rt, EXE_MEM_Rd, EXE_MEM_RegWrite, MEM_WB_Rd, MEM_WB_RegWrite, clk);
	// alu controlUnitd
	 
  
// EXE_MEM_Register
	EXE_MEM_Register exememr(EXE_MEM_Result, EXE_MEM_BranchAddress, EXE_MEM_DstReg, EXE_MEM_Rd, EXE_MEM_Zero, EXE_MEM_Rt, EXE_MEM_BranchEqual, EXE_MEM_BranchnotEqual,
								    EXE_MEM_MemRead, EXE_MEM_MemWrite, EXE_MEM_MemtoReg, EXE_MEM_RegWrite, EXE_BranchAddress, ALUOut_EXEC, EXE_DstReg, ID_EXE_Rd, ID_EXE_Rt,
								    EXE_Zero, ID_EXE_BranchEqual, ID_EXE_BranchnotEqual, ID_EXE_MemRead, ID_EXE_MemWrite, ID_EXE_MemtoReg, ID_EXE_RegWrite, clk);

// MEM Stage
	DataMemory DMem(MEM_Result, EXE_MEM_Result, EXE_MEM_Rt, EXE_MEM_MemRead, EXE_MEM_MemWrite, clk);
	BranchEqualAnd beand (BranchEqualResult, EXE_MEM_Zero, EXE_MEM_BranchEqual);
	BranchnotEqualAnd bneand(BranchnotEqualResult, EXE_MEM_Zero, EXE_MEM_BranchnotEqual);
	AddressOr addor (PC_Src, BranchEqualResult, BranchnotEqualResult);
	
// MEM_WB_Register
	MEM_WB_Register memwbreg (MEM_WB_MemData, MEM_WB_ALUData, MEM_WB_Rd, MEM_WB_DstReg, MEM_WB_MemtoReg, MEM_WB_RegWrite, MEM_Result, EXE_MEM_Result,
						           EXE_MEM_Rd, EXE_MEM_DstReg, EXE_MEM_MemtoReg, EXE_MEM_RegWrite, clk);
   	
// WB Stage
	WB_MUX wbmux (WB_Data, MEM_WB_MemData, MEM_WB_ALUData, MemtoReg, clk);
	
endmodule

module tst_2; 
	reg [31:0]PC_VALUE_;		  
	reg [31:0] cycle;
	Top top(PC_VALUE_);
	initial begin
		PC_VALUE_ <= 200;	  
		cycle <= 1;
	end				   
	always @(posedge top.clk) begin	

	if (cycle == 1)
	begin
		$display("cycle: %d" , cycle);
		$display("PC: %d",top.program_counter);				   
		$display("ALUOut_EXEC: %d" , top.ALUOut_EXEC);
		$display("$s1: %d" , top.regFile.registers_i[19], " The correct value is 5");
		$display("$s2: %d" , top.regFile.registers_i[20], " The correct value is 10");		
		$display("$s3: %d" , top.regFile.registers_i[21], " The correct value is 3");		
		$display("$s4: %d" , top.regFile.registers_i[22], " The correct value is 2");
		$display("$s5: %d" , top.regFile.registers_i[23], " The correct value is 15");
		$display("$s6: %d" , top.regFile.registers_i[24], " The correct value is -2  *** Check reporesentation");		
				
		
		end
			cycle = cycle + 1;
		
		
	end
endmodule
