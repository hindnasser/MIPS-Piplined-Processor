module Top (PC_value);

input PC_value;



endmodule
